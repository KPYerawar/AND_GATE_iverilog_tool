module gate (
    input A,
    input B,
    output Y
);
    and (Y, A, B);  // AND gate implementation
endmodule
